Analise de frequency response no V6
Vs   1    0   DC 0 AC 1 SIN(0 1 1000)
R1   1    2   1.02166163214k
R2   2    3   2.05713464724k 
R3   2    5   3.10288701080k 
R4   0    5   4.16870321182k 
R5   5    6   3.01167607597k 
R6   0   7.1  2.04520070018k 
Ve  7.1  7.2  0.00000000000  ;Fonte nula para medir a corrente
R7  7.2   8   1.02576029486k 

Cc   6    8   1.00334118042u ;Condensador C

Hd  5 8  Ve   8.29202733390k ;Fonte de voltagem
Gb  6 3 (2,5) 7.24529394385m ;Fonte de corrente


.ac DEC 100 0.1 1000000


.control
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

run
hardcopy plotmagnitude.ps db(V(6)) db(V(6)-V(8)) db(V(1))
hardcopy plotfase.ps 180/pi*ph(v(6)) 180/pi*ph(v(6)-v(8)) 180/pi*ph(v(1)) 

quit

.endc

.end

