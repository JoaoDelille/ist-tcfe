T4 Laboratory Simulation Results
.options savecurrents
.param Rin_value=100
.param Ci_value=365u
.param R1_value=80000
.param R2_value=20000
.param Rc_value=980
.param Re_value=1015
.param Cb_value=4390u
.param Rout_value=2335
.param Co_value=2250u
.param RL_value=8

.csparam Rin_value={Rin_value}
.csparam Ci_value={Ci_value}
.csparam R1_value={R1_value}
.csparam R2_value={R2_value}
.csparam Rc_value={Rc_value}
.csparam Re_value={Re_value}
.csparam Cb_value={Cb_value}
.csparam Rout_value={Rout_value}
.csparam Co_value={Co_value}
.csparam RL_value={RL_value}

.options savecurrents

* PHILIPS BJT'S
.MODEL BC557A PNP(IS=2.059E-14 ISE=2.971f    ISC=1.339E-14 XTI=3 BF=227.3 BR=7.690 IKF=0.08719 IKR=0.07646 XTB=1.5 VAF=37.2 VAR=11.42 VJE=0.5912 VJC=0.1 RE=0.6880 RC=0.6437 RB=1 RBM=1 IRB=1E-06 CJE=1.40E-11 CJC=1.113E-11 XCJC=0.6288 FC=0.7947 NF=1.003 NR=1.007 NE=1.316 NC=1.150 MJE=0.3572 MJC=0.3414 TF=7.046E-10 TR=1m2 ITF=0.1947 VTF=5.367 XTF=4.217 EG=1.11)
.MODEL BC547A NPN(IS=1.533E-14 ISE=7.932E-16 ISC=8.305E-14 XTI=3 BF=178.7 BR=8.628 IKF=0.12160 IKR=0.11210 XTB=1.5 VAF=69.7 VAR=44.70 VJE=0.4209 VJC=0.2 RE=0.6395 RC=0.6508 RB=1 RBM=1 IRB=1E-06 CJE=1.61E-11 CJC=4.388p    XCJC=0.6193 FC=0.7762 NF=1.002 NR=1.004 NE=1.436 NC=1.207 MJE=0.3071 MJC=0.2793 TF=4.995E-10 TR=1m2 ITF=0.7021 VTF=3.523 XTF=139.0 EG=1.11)

Vcc vcc 0 12.0
Vin in 0 0 ac 1.0 sin(0 10m 1k)
Rin in in2 {Rin_value}

* input coupling capacitor
Ci in2 base {Ci_value}

* bias circuit
R1 vcc base {R1_value}
R2 base 0 {R2_value}

* gain stage
Q1 coll base emit BC547A
Rc vcc coll {Rc_value}
Re emit 0 {Re_value}

* bypass capacitor
Cb emit 0 {Cb_value}

* output stage
Q2 0 coll emit2 BC557A
Rout emit2 vcc {Rout_value}

* output coupling capacitor
Co emit2 out {Co_value}

* load
RL out 0 8 {RL_value}

.op
.end

.control
set hcopypscolor=1
print all

* time analysis
tran 1e-5 1e-2
hardcopy vo1.ps vdb(coll)


* frequency analysis
ac dec 10 0.10 100MEG



hardcopy vo1f.ps vdb(coll)

hardcopy vo1f2.ps vp(coll)


hardcopy vo2f.ps vdb(out)

hardcopy vo2f2.ps vp(out)


let gain = db(v(out)[40]/v(in)[40])
hardcopy gain.ps db(v(out)/v(in))
hardcopy gain2.ps ph(v(out)/v(in))


meas AC wanted MAX vdb(out)
let ref=wanted-3

meas AC low WHEN vdb(out) = ref
meas AC up WHEN vdb(out) = ref CROSS=LAST


let resist=(Rin_value+R1_value+R2_value+Rc_value+Re_value+Rout_value+RL_value)*0.001
let capac=(Ci_value+Cb_value+Co_value)*1000000
let trans=2
let bandwidth=up-low
let cost=resist+capac+trans*0.1
let merit=((gain*bandwidth)/(cost*low))


echo "merit_TAB"
print low
print cost
print gain
print bandwidth
print merit
echo "merit_END"




let VCE=v(coll)-v(emit)
let VBE=v(base)-v(emit)
let VEB=v(emit2)-0
let VEC=v(emit2)-v(coll)

echo "op_TAB"
print VEC
print VEB
print VCE
print VBE
echo "op_END"



*input impedance in kohm
let Zin=abs(v(in2)[40]/vin#branch[40]/(-1000))

echo "input_TAB"
print Zin
echo "input_END"


quit
.endc
 
.end
