Final contender for the circuit, further testing required for fine tuning

.model Default D 
********************************
Vs 2 3 SIN( 0 12.7 50 )    ;                             
*********envelope detector     ;                        
*full bridge rectifier   ;     ;
D1  2  5  Default    ;   ;     ;
D2  0  2  Default    ;   ;     ;
D3  0  3  Default    ;   ;     ;
D4  3  5  Default    ;   ;     ;
**********************   ;     ;
*Rc    1 5 0              ;     ;
Ct    5 0 1.2u       ;     ;                      
**************************     ;            
*****voltage limiter           ;                 
.include stack.cir ;           ;             
*Rlim 5 4 0.00      ;           ;
Xlim1 5 6 inout20  ;           ;
Xlim2 6 7 inout20  ;           ;
Xlim3 7 8 inout20  ;           ;
Xlim4 8 9 inout10  ;           ;
Dlim5 9 0 Default  ;           ;    
********************           ;
.model Default D               ;
********************************
**********************************************
.measure tran Vavg  AVG v(5) from=155 to=155.2   ;
.measure tran Vmin  MIN v(5) from=155 to=155.2   ;
.measure tran Vmax  MAX v(5) from=155 to=155.2   ;
**********************************************
************************************************
.control                                       ;
set hcopypscolor=1                             ;
run                                            ;
                                               ;
tran 0.0002 155.2 155                            ;
hardcopy out.ps (v(5)) (v(2)-v(3))             ;
                                               ;
                           ;
hardcopy zoom.ps (v(5)-12)                     ;
                                               ;
quit                                           ;
.endc                                          ;
************************************************
.end

