Analise do V6 forcado
.options savecurrents
Vs   1    0   SIN(0 1 1000 0 0 0)
R1   1    2   1.02166163214k
R2   2    3   2.05713464724k 
R3   2    5   3.10288701080k 
R4   0    5   4.16870321182k 
R5   5    6   3.01167607597k 
R6   0   7.1  2.04520070018k 
Ve  7.1  7.2  0.00000000000  ;Fonte nula para medir a corrente
R7  7.2   8   1.02576029486k 

Cc   6    8   1.00334118042u ;Condensador C

Hd  5 8  Ve   8.29202733390m ;Fonte de voltagem
Gb  6 3 (2,5) 7.24529394385m ;Fonte de corrente


.ic v(6)=8.763595 v(8)=0     ;Condicao inicial do C
.tran 0.001ms 20ms uic

.control
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0
run
hardcopy plotfinal.ps    v(1) v(6) ;e suposto ser isto?
quit
.endc

.end

